`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    00:49:22 04/03/2024 
// Design Name: 
// Module Name:    halfSubtractor 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module halfSubtractor(
    input a,
    input b,
    output diff,
    output borrow
    );
	 
	 assign diff = a^b;
	 assign borrow = ~a&b;


endmodule
